`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2023/07/04 14:02:37
// Design Name: 
// Module Name: attention
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module attention(input clk, rst

    );
    
    reg [15:0] query[0:15][0:15];
    reg [15:0] key[0:15][0:15];
    //reg [15:0] value[0:3][0:3];
    
    reg [15:0] QK [0:15][0:15];
    
    integer i, j, k;
    
    reg [4:0] qk_address1, qk_address2;
    reg mat_mul;
    reg [15:0] m1_data,  m2_data, m3_data, m4_data;
    
    reg [3:0] state, state_2, state_3;
    
    parameter idle = 4'b0000;
    parameter matmul = 4'b0001;
    parameter scale = 4'b0010;
    parameter finish = 4'b0011;
    
    wire [15:0] mul_num, sum_num;
    
    reg [15:0] scale_dk = 16'b0011010000000000; //0.25
    
    reg clk_2hz;
    reg cnt;
    always@(posedge clk)begin
        if(rst)begin
            clk_2hz = 1;
            cnt = 0;
        end
        else
            if(cnt == 1)
                clk_2hz = ~clk_2hz;
            else 
                cnt = ~cnt;
    end
    
    
    always@(posedge clk_2hz)begin
         if(rst)begin
            for(i = 0; i < 16; i=i+1)begin
                for(j = 0; j < 16; j=j+1)begin
                    QK[i][j] = 16'b0;
                end
            end
            query[0][0] = 16'b0000000000000000; //0
            query[0][1] = 16'b0011110000000000; //1
            query[0][2] = 16'b0100000000000000; //2
            query[0][3] = 16'b0100001000000000; //3            
            query[0][4] = 16'b0100010000000000; //4
            query[0][5] = 16'b0100010100000000; //5
            query[0][6] = 16'b0100011000000000; //6
            query[0][7] = 16'b0100011100000000; //7
            query[0][8] = 16'b0100100000000000; //8
            query[0][9] = 16'b0100100010000000; //9
            query[0][10] = 16'b0100100100000000; //10
            query[0][11] = 16'b0100100110000000; //11
            query[0][12] = 16'b0100101000000000; //12
            query[0][13] = 16'b0100101010000000; //13
            query[0][14] = 16'b0100101100000000; //14
            query[0][15] = 16'b0100101110000000; //15
            
            query[1][15]  = 16'b0000000000000000; //0
            query[1][1]  = 16'b0011110000000000; //1
            query[1][2]  = 16'b0100000000000000; //2
            query[1][3]  = 16'b0100001000000000; //3            
            query[1][4]  = 16'b0100010000000000; //4
            query[1][5]  = 16'b0100010100000000; //5
            query[1][6]  = 16'b0100011000000000; //6
            query[1][7]  = 16'b0100011100000000; //7
            query[1][8]  = 16'b0100100000000000; //8
            query[1][9]  = 16'b0100100010000000; //9
            query[1][10] = 16'b0100100100000000; //10
            query[1][11] = 16'b0100100110000000; //11
            query[1][12] = 16'b0100101000000000; //12
            query[1][13] = 16'b0100101010000000; //13
            query[1][14] = 16'b0100101100000000; //14
            query[1][0] = 16'b0100101110000000; //15
            
            query[2][0]  = 16'b0000000000000000; //0
            query[2][14]  = 16'b0011110000000000; //1
            query[2][13]  = 16'b0100000000000000; //2
            query[2][3]  = 16'b0100001000000000; //3            
            query[2][4]  = 16'b0100010000000000; //4
            query[2][5]  = 16'b0100010100000000; //5
            query[2][6]  = 16'b0100011000000000; //6
            query[2][7]  = 16'b0100011100000000; //7
            query[2][8]  = 16'b0100100000000000; //8
            query[2][9]  = 16'b0100100010000000; //9
            query[2][10] = 16'b0100100100000000; //10
            query[2][11] = 16'b0100100110000000; //11
            query[2][12] = 16'b0100101000000000; //12
            query[2][2] = 16'b0100101010000000; //13
            query[2][1] = 16'b0100101100000000; //14
            query[2][15] = 16'b0100101110000000; //15
            
            query[3][0]  = 16'b0000000000000000; //0
            query[3][1]  = 16'b0011110000000000; //1
            query[3][2]  = 16'b0100000000000000; //2
            query[3][3]  = 16'b0100001000000000; //3            
            query[3][7]  = 16'b0100010000000000; //4
            query[3][6]  = 16'b0100010100000000; //5
            query[3][5]  = 16'b0100011000000000; //6
            query[3][4]  = 16'b0100011100000000; //7
            query[3][8]  = 16'b0100100000000000; //8
            query[3][9]  = 16'b0100100010000000; //9
            query[3][10] = 16'b0100100100000000; //10
            query[3][11] = 16'b0100100110000000; //11
            query[3][12] = 16'b0100101000000000; //12
            query[3][13] = 16'b0100101010000000; //13
            query[3][14] = 16'b0100101100000000; //14
            query[3][15] = 16'b0100101110000000; //15

            query[4][0]  = 16'b0100010000000000; 
            query[4][1]  = 16'b0100010100000000; 
            query[4][2]  = 16'b0100011000000000; 
            query[4][3]  = 16'b0100011100000000;           
            query[4][5]  = 16'b0100100000000000; 
            query[4][6]  = 16'b0100100010000000; 
            query[4][7]  = 16'b0100100100000000; 
            query[4][4]  = 16'b0100100110000000; 
            query[4][8]  = 16'b0100101000000000; 
            query[4][9]  = 16'b0100101010000000; 
            query[4][10] = 16'b0100101100000000; 
            query[4][11] = 16'b0100101110000000; 
            query[4][12] = 16'b0000000000000000; 
            query[4][13] = 16'b0011110000000000;
            query[4][14] = 16'b0100000000000000;
            query[4][15] = 16'b0100001000000000;
           
            query[5][2]  = 16'b0100010000000000; 
            query[5][3]  = 16'b0100010100000000; 
            query[5][0]  = 16'b0100011000000000; 
            query[5][1]  = 16'b0100011100000000;            
            query[5][4]  = 16'b0100100000000000; 
            query[5][5]  = 16'b0100100010000000; 
            query[5][6]  = 16'b0100100100000000; 
            query[5][7]  = 16'b0100100110000000; 
            query[5][8]  = 16'b0100101000000000; 
            query[5][9]  = 16'b0100101010000000; 
            query[5][10] = 16'b0100101100000000; 
            query[5][11] = 16'b0100101110000000; 
            query[5][12] = 16'b0000000000000000; 
            query[5][13] = 16'b0011110000000000; 
            query[5][14] = 16'b0100000000000000; 
            query[5][15] = 16'b0100001000000000; 
          
            query[6][0]  = 16'b0100010000000000; 
            query[6][1]  = 16'b0100010100000000; 
            query[6][2]  = 16'b0100011000000000; 
            query[6][3]  = 16'b0100011100000000;            
            query[6][4]  = 16'b0100100000000000; 
            query[6][5]  = 16'b0100100010000000; 
            query[6][6]  = 16'b0100100100000000; 
            query[6][7]  = 16'b0100100110000000; 
            query[6][8]  = 16'b0100101000000000; 
            query[6][9]  = 16'b0100101010000000; 
            query[6][10] = 16'b0100101100000000; 
            query[6][11] = 16'b0100101110000000; 
            query[6][12] = 16'b0000000000000000; 
            query[6][13] = 16'b0011110000000000; 
            query[6][14] = 16'b0100000000000000; 
            query[6][15] = 16'b0100001000000000; 
          
            query[7][0]  = 16'b0100010000000000; 
            query[7][1]  = 16'b0100010100000000; 
            query[7][2]  = 16'b0100011000000000; 
            query[7][3]  = 16'b0100011100000000;            
            query[7][4]  = 16'b0100100000000000; 
            query[7][5]  = 16'b0100100010000000; 
            query[7][6]  = 16'b0100100100000000; 
            query[7][7]  = 16'b0100100110000000; 
            query[7][8]  = 16'b0100101000000000; 
            query[7][9]  = 16'b0100101010000000; 
            query[7][10] = 16'b0100101100000000; 
            query[7][11] = 16'b0100101110000000; 
            query[7][12] = 16'b0000000000000000; 
            query[7][13] = 16'b0011110000000000; 
            query[7][15] = 16'b0100000000000000; 
            query[7][14] = 16'b0100001000000000; 
            
            query[8][0]  = 16'b0100100010000000; //0
            query[8][1]  = 16'b0100100100000000; //1
            query[8][2]  = 16'b0100100110000000; //2
            query[8][3]  = 16'b0100101000000000; //3            
            query[8][4]  = 16'b0100101010000000; //4
            query[8][5]  = 16'b0100101100000000; //5
            query[8][6]  = 16'b0100101110000000; //6
            query[8][7]  = 16'b0000000000000000; //7
            query[8][8]  = 16'b0011110000000000; //8
            query[8][9]  = 16'b0100000000000000; //9
            query[8][10] = 16'b0100001000000000; //10
            query[8][11] = 16'b0100010000000000; //11
            query[8][13] = 16'b0100010100000000; //12
            query[8][14] = 16'b0100011000000000; //13
            query[8][15] = 16'b0100011100000000; //14
            query[8][12] = 16'b0100100000000000; //15
            
            query[9][0]  = 16'b0100100010000000; //0
            query[9][2]  = 16'b0100100100000000; //1
            query[9][3]  = 16'b0100100110000000; //2
            query[9][1]  = 16'b0100101000000000; //3            
            query[9][4]  = 16'b0100101010000000; //4
            query[9][5]  = 16'b0100101100000000; //5
            query[9][6]  = 16'b0100101110000000; //6
            query[9][7]  = 16'b0000000000000000; //7
            query[9][8]  = 16'b0011110000000000; //8
            query[9][9]  = 16'b0100000000000000; //9
            query[9][10] = 16'b0100001000000000; //10
            query[9][11] = 16'b0100010000000000; //11
            query[9][12] = 16'b0100010100000000; //12
            query[9][13] = 16'b0100011000000000; //13
            query[9][14] = 16'b0100011100000000; //14
            query[9][15] = 16'b0100100000000000; //15
            
            query[10][0]  = 16'b0100100010000000; //0
            query[10][1]  = 16'b0100100100000000; //1
            query[10][2]  = 16'b0100100110000000; //2
            query[10][4]  = 16'b0100101000000000; //3            
            query[10][3]  = 16'b0100101010000000; //4
            query[10][5]  = 16'b0100101100000000; //5
            query[10][6]  = 16'b0100101110000000; //6
            query[10][7]  = 16'b0000000000000000; //7
            query[10][8]  = 16'b0011110000000000; //8
            query[10][9]  = 16'b0100000000000000; //9
            query[10][10] = 16'b0100001000000000; //10
            query[10][11] = 16'b0100010000000000; //11
            query[10][12] = 16'b0100010100000000; //12
            query[10][13] = 16'b0100011000000000; //13
            query[10][14] = 16'b0100011100000000; //14
            query[10][15] = 16'b0100100000000000; //15
            
            query[11][0]  = 16'b0100100010000000; //0
            query[11][1]  = 16'b0100100100000000; //1
            query[11][2]  = 16'b0100100110000000; //2
            query[11][3]  = 16'b0100101000000000; //3            
            query[11][4]  = 16'b0100101010000000; //4
            query[11][5]  = 16'b0100101100000000; //5
            query[11][6]  = 16'b0100101110000000; //6
            query[11][7]  = 16'b0000000000000000; //7
            query[11][8]  = 16'b0011110000000000; //8
            query[11][9]  = 16'b0100000000000000; //9
            query[11][10] = 16'b0100001000000000; //10
            query[11][11] = 16'b0100010000000000; //11
            query[11][12] = 16'b0100010100000000; //12
            query[11][13] = 16'b0100011000000000; //13
            query[11][14] = 16'b0100011100000000; //14
            query[11][15] = 16'b0100100000000000; //15
            
            query[12][1]  = 16'b0100101000000000; //0
            query[12][2]  = 16'b0100101010000000; //1
            query[12][0]  = 16'b0100101100000000; //2
            query[12][3]  = 16'b0100101110000000; //3            
            query[12][4]  = 16'b0000000000000000; //4
            query[12][5]  = 16'b0011110000000000; //5
            query[12][6]  = 16'b0100000000000000; //6
            query[12][7]  = 16'b0100001000000000; //7
            query[12][8]  = 16'b0100010000000000; //8
            query[12][9]  = 16'b0100010100000000; //9
            query[12][10] = 16'b0100011000000000; //10
            query[12][11] = 16'b0100011100000000; //11
            query[12][12] = 16'b0100100000000000; //
            query[12][13] = 16'b0100100010000000; //
            query[12][14] = 16'b0100100100000000; //
            query[12][15] = 16'b0100100110000000; //
            
            query[13][0]  = 16'b0100101000000000; //0
            query[13][1]  = 16'b0100101010000000; //1
            query[13][2]  = 16'b0100101100000000; //2
            query[13][5]  = 16'b0100101110000000; //3            
            query[13][4]  = 16'b0000000000000000; //4
            query[13][3]  = 16'b0011110000000000; //5
            query[13][6]  = 16'b0100000000000000; //6
            query[13][7]  = 16'b0100001000000000; //7
            query[13][8]  = 16'b0100010000000000; //8
            query[13][9]  = 16'b0100010100000000; //9
            query[13][10] = 16'b0100011000000000; //10
            query[13][11] = 16'b0100011100000000; //11
            query[13][12] = 16'b0100100000000000; //12
            query[13][13] = 16'b0100100010000000; //13
            query[13][14] = 16'b0100100100000000; //14
            query[13][15] = 16'b0100100110000000; //15
            
            query[14][0]  = 16'b0100101000000000; //0
            query[14][1]  = 16'b0100101010000000; //1
            query[14][2]  = 16'b0100101100000000; //2
            query[14][3]  = 16'b0100101110000000; //3            
            query[14][4]  = 16'b0000000000000000; //4
            query[14][5]  = 16'b0011110000000000; //5
            query[14][6]  = 16'b0100000000000000; //6
            query[14][7]  = 16'b0100001000000000; //7
            query[14][8]  = 16'b0100010000000000; //8
            query[14][9]  = 16'b0100010100000000; //9
            query[14][10] = 16'b0100011000000000; //10
            query[14][11] = 16'b0100011100000000; //11
            query[14][12] = 16'b0100100000000000; //12
            query[14][13] = 16'b0100100010000000; //13
            query[14][15] = 16'b0100100100000000; //14
            query[14][14] = 16'b0100100110000000; //15
            
            query[15][0]  = 16'b0100101000000000; //0
            query[15][1]  = 16'b0100101010000000; //1
            query[15][2]  = 16'b0100101100000000; //2
            query[15][3]  = 16'b0100101110000000; //3            
            query[15][4]  = 16'b0000000000000000; //4
            query[15][5]  = 16'b0011110000000000; //5
            query[15][6]  = 16'b0100000000000000; //6
            query[15][7]  = 16'b0100001000000000; //7
            query[15][8]  = 16'b0100010000000000; //8
            query[15][9]  = 16'b0100010100000000; //9
            query[15][10] = 16'b0100011000000000; //10
            query[15][11] = 16'b0100011100000000; //11
            query[15][12] = 16'b0100100000000000; //12
            query[15][13] = 16'b0100100010000000; //13
            query[15][14] = 16'b0100100100000000; //14
            query[15][15] = 16'b0100100110000000; //15
            
            key[0][0] =   16'b0010111001100110; //0.1
            key[0][1] =   16'b0011001001100110; //0.2
            key[0][2] =   16'b0011010011001101; //0.3
            key[0][3] =   16'b0011011001100110; //0.4
            key[0][4] =   16'b0011100000000000; //0.5
            key[0][5] =   16'b0011100011001101; //0.6
            key[0][6] =   16'b0011100110011010; //0.7
            key[0][7] =   16'b0011101001100110; //0.8
            key[0][8] =   16'b0011101100110011; //0.9
            key[0][9] =   16'b1010111100001010; //-0.11
            key[0][10] =  16'b1010111110101110; //-0.12
            key[0][11] =  16'b1011000000101001; //-0.13
            key[0][12] =  16'b1011000001111011; //-0.14
            key[0][13] =  16'b1011000011001101; //-0.15
            key[0][14] =  16'b1011000011001101; //-0.15
            key[0][15] =  16'b1011000011001101; //-0.15
            
            key[1][0]  =  16'b0010111100001010; //0.1
            key[1][1]  =  16'b0011001010111000; //0.2
            key[1][2]  =  16'b0011010011110110; //0.3
            key[1][3]  =  16'b0011011010001111; //0.4
            key[1][4]  =  16'b0011100000010100; //0.5
            key[1][5]  =  16'b0011100011100001; //0.6
            key[1][6]  =  16'b0011100110101110; //0.7
            key[1][7]  =  16'b0011101001111011; //0.8
            key[1][8]  =  16'b0011101101000111; //0.9
            key[1][9]  =  16'b1010111100011010; //-0.11
            key[1][10] =  16'b1010111110111110; //-0.12
            key[1][11] =  16'b1011000000110001; //-0.13
            key[1][12] =  16'b1011000010000011; //-0.14
            key[1][13] =  16'b1011000011010101; //-0.15
            key[1][14] =  16'b1011000011010101; //-0.15
            key[1][15] =  16'b1011000011010101; //-0.15
            
            key[2][0]  =  16'b0011110001100110; //0.1
            key[2][1]  =  16'b0100000001100110; //0.2
            key[2][2]  =  16'b0100001010011010; //0.3
            key[2][3]  =  16'b0100010001100110; //0.4
            key[2][4]  =  16'b0100010110000000; //0.5
            key[2][5]  =  16'b0100011010011010; //0.6
            key[2][6]  =  16'b0100011110110011; //0.7
            key[2][7]  =  16'b0100100001100110; //0.8
            key[2][8]  =  16'b0100100011110011; //0.9
            key[2][9]  =  16'b1100100100001110; //-0.11
            key[2][10] =  16'b1100100100001111; //-0.12
            key[2][11] =  16'b1100100100010000; //-0.13
            key[2][12] =  16'b1100100100010010; //-0.14
            key[2][13] =  16'b1100100100010011; //-0.15
            key[2][14] =  16'b1100100100010011; //-0.15
            key[2][15] =  16'b1100100100010011; //-0.15
            
            key[3][0]  =  16'b0100110100000110; 
            key[3][1]  =  16'b0100110100001101; 
            key[3][2]  =  16'b0100110100010011; 
            key[3][3]  =  16'b0100110100011010; 
            key[3][4]  =  16'b0100110100100000; 
            key[3][5]  =  16'b0100110100100110; 
            key[3][6]  =  16'b0100110100101101; 
            key[3][7]  =  16'b0100110100110011; 
            key[3][8]  =  16'b0100110100111010; 
            key[3][9]  =  16'b1100110100000111; 
            key[3][10] =  16'b1100110100000111; 
            key[3][11] =  16'b1100110100001000; 
            key[3][12] =  16'b1100110100001001; 
            key[3][13] =  16'b1100110100001010; 
            key[3][14] =  16'b1100110100001010; 
            key[3][15] =  16'b1100110100001010; 
           
            key[4][1]  =  16'b0010111001100110; 
            key[4][0]  =  16'b0011001001100110; 
            key[4][2]  =  16'b0011010011001101; 
            key[4][3]  =  16'b0011011001100110; 
            key[4][4]  =  16'b0011100000000000; 
            key[4][5]  =  16'b0011100011001101; 
            key[4][6]  =  16'b0011100110011010; 
            key[4][7]  =  16'b0011101001100110; 
            key[4][8]  =  16'b0011101100110011; 
            key[4][9]  =  16'b1010111100001010; 
            key[4][10] =  16'b1010111110101110; 
            key[4][11] =  16'b1011000000101001; 
            key[4][12] =  16'b1011000001111011; 
            key[4][13] =  16'b1011000011001101; 
            key[4][14] =  16'b1011000011001101; 
            key[4][15] =  16'b1011000011001101; 
           
            key[5][1]  =  16'b0010111100001010; 
            key[5][0]  =  16'b0011001010111000; 
            key[5][2]  =  16'b0011010011110110; 
            key[5][3]  =  16'b0011011010001111; 
            key[5][4]  =  16'b0011100000010100; 
            key[5][5]  =  16'b0011100011100001; 
            key[5][6]  =  16'b0011100110101110; 
            key[5][7]  =  16'b0011101001111011; 
            key[5][8]  =  16'b0011101101000111; 
            key[5][9]  =  16'b1010111100011010; 
            key[5][10] =  16'b1010111110111110; 
            key[5][11] =  16'b1011000000110001; 
            key[5][12] =  16'b1011000010000011; 
            key[5][13] =  16'b1011000011010101; 
            key[5][14] =  16'b1011000011010101; 
            key[5][15] =  16'b1011000011010101; 
           
            key[6][1]  =  16'b0011110001100110; 
            key[6][0]  =  16'b0100000001100110; 
            key[6][2]  =  16'b0100001010011010; 
            key[6][3]  =  16'b0100010001100110; 
            key[6][4]  =  16'b0100010110000000; 
            key[6][5]  =  16'b0100011010011010; 
            key[6][6]  =  16'b0100011110110011; 
            key[6][7]  =  16'b0100100001100110; 
            key[6][8]  =  16'b0100100011110011; 
            key[6][9]  =  16'b1100100100001110; 
            key[6][10] =  16'b1100100100001111; 
            key[6][11] =  16'b1100100100010000; 
            key[6][12] =  16'b1100100100010010; 
            key[6][13] =  16'b1100100100010011; 
            key[6][14] =  16'b1100100100010011; 
            key[6][15] =  16'b1100100100010011; 
           
            key[7][1]  =  16'b0100110100000110; 
            key[7][0]  =  16'b0100110100001101; 
            key[7][2]  =  16'b0100110100010011; 
            key[7][3]  =  16'b0100110100011010; 
            key[7][4]  =  16'b0100110100100000; 
            key[7][5]  =  16'b0100110100100110; 
            key[7][6]  =  16'b0100110100101101; 
            key[7][7]  =  16'b0100110100110011; 
            key[7][8]  =  16'b0100110100111010; 
            key[7][9]  =  16'b1100110100000111; 
            key[7][10] =  16'b1100110100000111; 
            key[7][11] =  16'b1100110100001000; 
            key[7][12] =  16'b1100110100001001; 
            key[7][13] =  16'b1100110100001010; 
            key[7][14] =  16'b1100110100001010; 
            key[7][15] =  16'b1100110100001010; 
            
            key[8][0]  =  16'b0010111001100110;
            key[8][1]  =  16'b0011001001100110;
            key[8][3]  =  16'b0011010011001101;
            key[8][2]  =  16'b0011011001100110;
            key[8][4]  =  16'b0011100000000000;
            key[8][5]  =  16'b0011100011001101;
            key[8][6]  =  16'b0011100110011010;
            key[8][7]  =  16'b0011101001100110;
            key[8][8]  =  16'b0011101100110011;
            key[8][9]  =  16'b1010111100001010;
            key[8][10] =  16'b1010111110101110;
            key[8][11] =  16'b1011000000101001;
            key[8][12] =  16'b1011000001111011;
            key[8][13] =  16'b1011000011001101;
            key[8][14] =  16'b1011000011001101;
            key[8][15] =  16'b1011000011001101;
                                              
            key[9][0]  =  16'b0010111100001010;
            key[9][1]  =  16'b0011001010111000;
            key[9][3]  =  16'b0011010011110110;
            key[9][2]  =  16'b0011011010001111;
            key[9][4]  =  16'b0011100000010100;
            key[9][5]  =  16'b0011100011100001;
            key[9][6]  =  16'b0011100110101110;
            key[9][7]  =  16'b0011101001111011;
            key[9][8]  =  16'b0011101101000111;
            key[9][9]  =  16'b1010111100011010;
            key[9][10] =  16'b1010111110111110;
            key[9][11] =  16'b1011000000110001;
            key[9][12] =  16'b1011000010000011;
            key[9][13] =  16'b1011000011010101;
            key[9][14] =  16'b1011000011010101;
            key[9][15] =  16'b1011000011010101;
                                              
            key[10][0]  = 16'b0011110001100110;
            key[10][1]  = 16'b0100000001100110;
            key[10][3]  = 16'b0100001010011010;
            key[10][2]  = 16'b0100010001100110;
            key[10][4]  = 16'b0100010110000000;
            key[10][5]  = 16'b0100011010011010;
            key[10][6]  = 16'b0100011110110011;
            key[10][7]  = 16'b0100100001100110;
            key[10][8]  = 16'b0100100011110011;
            key[10][9]  = 16'b1100100100001110;
            key[10][10] = 16'b1100100100001111;
            key[10][11] = 16'b1100100100010000;
            key[10][12] = 16'b1100100100010010;
            key[10][13] = 16'b1100100100010011;
            key[10][14] = 16'b1100100100010011;
            key[10][15] = 16'b1100100100010011;
                                              
            key[11][0]  = 16'b0100110100000110;
            key[11][1]  = 16'b0100110100001101;
            key[11][3]  = 16'b0100110100010011;
            key[11][2]  = 16'b0100110100011010;
            key[11][4]  = 16'b0100110100100000;
            key[11][5]  = 16'b0100110100100110;
            key[11][6]  = 16'b0100110100101101;
            key[11][7]  = 16'b0100110100110011;
            key[11][8]  = 16'b0100110100111010;
            key[11][9]  = 16'b1100110100000111;
            key[11][10] = 16'b1100110100000111;
            key[11][11] = 16'b1100110100001000;
            key[11][12] = 16'b1100110100001001;
            key[11][13] = 16'b1100110100001010;
            key[11][14] = 16'b1100110100001010;
            key[11][15] = 16'b1100110100001010;
                                              
            key[12][0]  = 16'b0010111001100110;
            key[12][1]  = 16'b0011001001100110;
            key[12][2]  = 16'b0011010011001101;
            key[12][3]  = 16'b0011011001100110;
            key[12][5]  = 16'b0011100000000000;
            key[12][4]  = 16'b0011100011001101;
            key[12][6]  = 16'b0011100110011010;
            key[12][7]  = 16'b0011101001100110;
            key[12][8]  = 16'b0011101100110011;
            key[12][9]  = 16'b1010111100001010;
            key[12][10] = 16'b1010111110101110;
            key[12][11] = 16'b1011000000101001;
            key[12][12] = 16'b1011000001111011;
            key[12][13] = 16'b1011000011001101;
            key[12][14] = 16'b1011000011001101;
            key[12][15] = 16'b1011000011001101;
                                              
            key[13][0]  = 16'b0010111100001010;
            key[13][1]  = 16'b0011001010111000;
            key[13][2]  = 16'b0011010011110110;
            key[13][3]  = 16'b0011011010001111;
            key[13][5]  = 16'b0011100000010100;
            key[13][4]  = 16'b0011100011100001;
            key[13][6]  = 16'b0011100110101110;
            key[13][7]  = 16'b0011101001111011;
            key[13][8]  = 16'b0011101101000111;
            key[13][9]  = 16'b1010111100011010;
            key[13][10] = 16'b1010111110111110;
            key[13][11] = 16'b1011000000110001;
            key[13][12] = 16'b1011000010000011;
            key[13][13] = 16'b1011000011010101;
            key[13][14] = 16'b1011000011010101;
            key[13][15] = 16'b1011000011010101;
                                              
            key[14][0]  = 16'b0011110001100110;
            key[14][1]  = 16'b0100000001100110;
            key[14][2]  = 16'b0100001010011010;
            key[14][3]  = 16'b0100010001100110;
            key[14][5]  = 16'b0100010110000000;
            key[14][4]  = 16'b0100011010011010;
            key[14][6]  = 16'b0100011110110011;
            key[14][7]  = 16'b0100100001100110;
            key[14][8]  = 16'b0100100011110011;
            key[14][9]  = 16'b1100100100001110;
            key[14][10] = 16'b1100100100001111;
            key[14][11] = 16'b1100100100010000;
            key[14][12] = 16'b1100100100010010;
            key[14][13] = 16'b1100100100010011;
            key[14][14] = 16'b1100100100010011;
            key[14][15] = 16'b1100100100010011;
                                              
            key[15][0]  = 16'b0100110100000110;
            key[15][1]  = 16'b0100110100001101;
            key[15][2]  = 16'b0100110100010011;
            key[15][3]  = 16'b0100110100011010;
            key[15][5]  = 16'b0100110100100000;
            key[15][4]  = 16'b0100110100100110;
            key[15][6]  = 16'b0100110100101101;
            key[15][7]  = 16'b0100110100110011;
            key[15][8]  = 16'b0100110100111010;
            key[15][9]  = 16'b1100110100000111;
            key[15][10] = 16'b1100110100000111;
            key[15][11] = 16'b1100110100001000;
            key[15][12] = 16'b1100110100001001;
            key[15][13] = 16'b1100110100001010;
            key[15][14] = 16'b1100110100001010;
            key[15][15] = 16'b1100110100001010;
            
            m1_data = 16'b0;
            m2_data = 16'b0;
            m3_data = 16'b0;
            m4_data = 16'b0;
            i = 0;
            j = 0;
            k = 0;
            mat_mul = 0;
            state <= 4'b1;
            state_2 <= 4'b0;
            state_3 <= 4'b0;
         end
         else begin
         case(state) 
            4'b0001:begin
                case(state_2)
                    2'b00: begin
                        if( k < 16) begin
                            if(j < 16) begin
                                qk_address1 = i;
                                qk_address2 = k;
                                m1_data = query[i][j];
                                m2_data = key[k][j];                                   
                                state_2 = 1;
                            end
                            else begin
                                j = 0;
                                k = k + 1;
                            end
                        end
                        else begin
                            i = i + 1;
                            j = 0;
                            k = 0;
                            if(i == 16)begin
                                i = 0;
                                state = state + 1;
                            end
                        end
                    end
                    2'b01: begin
                            m3_data = QK[qk_address1][qk_address2];
                            m4_data = mul_num; 
                            state_2 = 2;
                    end
                    2'b10:begin
                        state_2 = 3;
                    end
                    2'b11:begin
                        QK[qk_address1][qk_address2] = sum_num;
                        j = j + 1;
                        state_2 = 0;
                    end
                endcase
            end
            4'b0010:begin
                case(state_3)
                    2'b00: begin
                        if(i < 16)
                            if(k < 16) begin
                                m1_data = QK[i][k];
                                m2_data = scale_dk;
                                state_3 = 1;
                            end
                            else begin
                                i = i + 1;
                                k = 0;
                            end
                        else begin
                            i = 0;
                            state = state + 1;
                        end
                    end
                    2'b01: begin
                        QK[i][k] = mul_num;
                        state_3 = 0;
                        k = k + 1;
                    end
                endcase
            end
         endcase
        end
    end
    
    /*
    matrix_multiplier mp(
    .clk(clk),
    .rst(rst),
    .mat_mul(mat_mul),
    .m1_address1(m1_address1),
    .m1_address2(m1_address2),
    .m1_data(m1_data),
    .m2_address1(m2_address1),
    .m2_address2(m2_address2),
    .m2_data(m2_data),
    .out_data()
    );*/
    
    signed_floating_point_multiplier SFPM(
    .operand_a(m1_data),
    .operand_b(m2_data),
    .clk(clk),
    .rst(rst),
    .result(mul_num)
);
    signed_floating_point_adder SFPA(
    .operand_a(m3_data),
    .operand_b(m4_data),
    .clk(clk),
    .rst(rst),
    .result(sum_num)
);
endmodule


